library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;

entity CharacterROM is
	port (
		i_Char		: in	std_logic_vector (7 downto 0);
		i_Clk		: in	std_logic;
		
		o_Dots		: out	std_logic_vector (95 downto 0)
	);
end CharacterROM;

architecture Behavioral of CharacterROM is
	type rom_type is array (95 downto 0) of std_logic_vector(49 downto 0);
	constant character_table : rom_type := (
		-- space
		"00000000000000000000000000000000000000000000000000",
		-- !
		"00100001000010000100001000000000100001000000000000",
		-- "
		"01010010100101000000000000000000000000000000000000",
		-- #
		"01010010101111101010111110101001010000000000000000",
		-- $
		"00100011111010001110001011111000100000000000000000",
		-- %
		"00000110011101000100010111001100000000000000000000",
		-- &
		"01100100101010001000101011001001101000000000000000",
		-- '
		"00100001000100000000000000000000000000000000000000",
		-- (
		"00010001000100001000010000010000010000000000000000",
		-- )
		"01000001000001000010000100010001000000000000000000",
		-- *
		"00000001001010101110101010010000000000000000000000",
		-- +
		"00000001000010011111001000010000000000000000000000",
		-- ,
		"00000000000000000000000000010000100010000000000000",
		-- -
		"00000000000000011111000000000000000000000000000000",
		-- .
		"00000000000000000000000000000000100001000000000000",
		-- /
		"00001000100001000100010000100010000000000000000000",
		-- 0
		"01110100011001110101110011000101110000000000000000",
		-- 1
		"00100011000010000100001000010001110000000000000000",
		-- 2
		"01110100010000100010001000100011111000000000000000",
		-- 3
		"01110100010000101110000011000101110000000000000000",
		-- 4
		"00010001100101010010111110001000111000000000000000",
		-- 5
		"11111100001111000001000011000101110000000000000000",
		-- 6
		"00110010001000011110100011000101110000000000000000",
		-- 7
		"11111000010001000100010000100001000000000000000000",
		-- 8
		"01110100011000101110100011000101110000000000000000",
		-- 9
		"01110100011000101111000010001001100000000000000000",
		-- :
		"00000001000010000000001000010000000000000000000000",
		-- ;
		"00000001000010000000001000010001000000000000000000",
		-- <
		"00010001000100010000010000010000010000000000000000",
		-- =
		"00000000001111100000111110000000000000000000000000",
		-- >
		"01000001000001000001000100010001000000000000000000",
		-- ?
		"01110100010000100010001000000000100000000000000000",
		-- @
		"01110100011001110101101011000001110000000000000000",
		-- A
		"01110100011000110001111111000110001000000000000000",
		-- B
		"11110100011000111110100011000111110000000000000000",
		-- C
		"01110100011000010000100001000101110000000000000000",
		-- D
		"11110100011000110001100011000111110000000000000000",
		-- E
		"11111100001000011110100001000011111000000000000000",
		-- F
		"11111100001000011110100001000010000000000000000000",
		-- G
		"01110100011000010011100011000101110000000000000000",
		-- H
		"10001100011000111111100011000110001000000000000000",
		-- I
		"01110001000010000100001000010001110000000000000000",
		-- J
		"11111000010000100001100011000101110000000000000000",
		-- K
		"10001100101010011000101001001010001000000000000000",
		-- L
		"10000100001000010000100001000011111000000000000000",
		-- M
		"10001110111010110101100011000110001000000000000000",
		-- N
		"10001100011100110101100111000110001000000000000000",
		-- O
		"01110100011000110001100011000101110000000000000000",
		-- P
		"11110100011000111110100001000010000000000000000000",
		-- Q
		"01110100011000110001101011001001101000000000000000",
		-- R
		"11110100011000111110101001001010001000000000000000",
		-- S
		"01110100011000001110000011000101110000000000000000",
		-- T
		"11111001000010000100001000010000100000000000000000",
		-- U
		"10001100011000110001100011000101110000000000000000",
		-- V
		"10001100011000110001100010101000100000000000000000",
		-- W
		"10001100011000110101101011101110001000000000000000",
		-- X
		"10001100010101000100010101000110001000000000000000",
		-- Y
		"10001100010101000100001000010000100000000000000000",
		-- Z
		"11111000010001000100010001000011111000000000000000",
		-- [
		"01110010000100001000010000100001110000000000000000",
		-- -Y-
		"10001010101111100100111110010000100000000000000000",
		-- ]
		"01110000100001000010000100001001110000000000000000",
		-- ^
		"00100010101000100000000000000000000000000000000000",
		-- _
		"00000000000000000000000000000011111000000000000000",
		-- `
		"01000001000001000000000000000000000000000000000000",
		-- a
		"00000000000111000001011111000101111000000000000000",
		-- b
		"10000100001011011001100011000111110000000000000000",
		-- c
		"00000000000111010001100001000101110000000000000000",
		-- d
		"00001000010110110011100011000101111000000000000000",
		-- e
		"00000000000111010001111111000001110000000000000000",
		-- f
		"00110010010100011100010000100001000000000000000000",
		-- g
		"00000000000111110001100010111100001111100000000000",
		-- h
		"10000100001011011001100011000110001000000000000000",
		-- i
		"00100000000110000100001000010001110000000000000000",
		-- j
		"00010000000001000010000100001010010011000000000000",
		-- k
		"10000100001001010100110001010010010000000000000000",
		-- l
		"01100001000010000100001000010001110000000000000000",
		-- m
		"00000000001101010101101011000110001000000000000000",
		-- n
		"00000000001011011001100011000110001000000000000000",
		-- o
		"00000000000111010001100011000101110000000000000000",
		-- p
		"00000000001111010001111101000010000000000000000000",
		-- q
		"00000000000110110011011110000100001000000000000000",
		-- r
		"00000000001011011001100001000010000000000000000000",
		-- s
		"00000000000111010000011100000111110000000000000000",
		-- t
		"01000010001111001000010000100100110000000000000000",
		-- u
		"00000000001000110001100011001101101000000000000000",
		-- v
		"00000000001000110001100010101000100000000000000000",
		-- w
		"00000000001000110001101011010101010000000000000000",
		-- x
		"00000000001000101010001000101010001000000000000000",
		-- y
		"00000000001000110001011110000111110000000000000000",
		-- z
		"00000000001111100010001000100011111000000000000000",
		-- {
		"00010001000010001000001000010000010000000000000000",
		-- |
		"00100001000010000100001000010000100000000000000000",
		-- }
		"01000001000010000010001000010001000000000000000000",
		-- ->
		"00000001000001011111000100010000000000000000000000",
		-- <-
		"00000001000100011111010000010000000000000000000000"
	);
	
	signal tmp_rd : std_logic_vector (49 downto 0);
begin
	
	-- Char data is 	5x10
	-- Output data is	8x12
	
	process (i_CLK)
	begin
		if rising_edge(i_CLK) then
			tmp_rd <= character_table(to_integer(unsigned(i_Char)) - 32);
		end if;
	end process;
	
	GEN_PADDING: for i in 0 to 9 generate
		o_Dots((i * 8 + 7) downto (i * 8)) <=
			tmp_rd((i * 5 + 4) downto (i * 5)) & "000";
	end generate GEN_PADDING;
	
	o_Dots(95 downto 80) <= (others => '0');
	
end Behavioral;
